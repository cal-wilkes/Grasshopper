library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lookup is
	port (  clk: in std_logic;
			reset: in std_logic;
			ones: in integer;
			tens: in integer;
			tenths: in integer;
			scan_line_x: in std_logic_vector(10 downto 0);
			scan_line_y: in std_logic_vector(10 downto 0);
			colour: in std_logic_vector(11 downto 0);
			tablevalue: in std_logic_vector(8 downto 0);
			red: out std_logic_vector(3 downto 0);
			blue: out std_logic_vector(3 downto 0);
			green: out std_logic_vector(3 downto 0)
			);
end lookup;


architecture behaviour of lookup is

type vec is array (13 downto 0) of std_logic;
type matrix is array(17 downto 0) of vec;

signal pixel_colour: std_logic_vector(11 downto 0);

signal i_ones: matrix;
signal i_tens: matrix;
signal i_tenths: matrix;

constant size: std_logic_vector:= "1000";
signal counter: std_logic_vector := size;				   
							   							
							   
constant nine: matrix:= 	   (
							   ('0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0','0','0'),	
							   ('0','0','0','0','1','1','1','1','1,1,1,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
							   (0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0)
							   );
							   
constant eight: matrix:= 		(
								(0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),	
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0)
								);
								
constant seven: matrix:= 		(
								(0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),		
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,1,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0)
								);
								
constant six: matrix:= 		  (
							  (0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),	
							  (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0)
							  );
							  
constant five: matrix:= 	   (
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),		
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
							   (0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0)
							   );
							   
constant four: matrix:= 	   (
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),	
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,1,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,1,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
							   (0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
							   (0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0)
							    );	
							   
constant three: matrix:= 		(
								(0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),	
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							    (0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0)
								);	
								
constant two: matrix:= 		  (
							  (0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0),	
							  (0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0),
							  (0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0),
							  (0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0)
							   );	
							  
constant one: matrix:= 		  (
							  (0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),		
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
							  (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0)
							   );
							  
constant zero: matrix:= 	   (
							   (0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0),		
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0,0,0),
							   (0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
							   (0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0)
							   );							   
						
							   
process: pixel(scan_line_x, scan_line_y)

							if(counter <= 1)then
								counter <= size;
							else
								pixel_colour <= colour when ((scan_line_x >= box_loc_x) and (scan_line_x < box_loc_x + box_width) and
															(scan_line_y >= box_loc_y) and (scan_line_y < box_loc_y + box_width)
							else
								pixel_colour <= "111111111111";
								
end process;

red <= pixel_colour(11 downto 8);
green <= pixel_colour(7 downto 4);
blue <= pixel_colour(3 downto 0);

end behaviour;
